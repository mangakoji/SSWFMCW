// SIN_TBL_s11_s11.v
//
//
//170522su      :debug C_XCLIP_1POINT0
//170516tu      :add EN_CK_i , CK&XARST add tail suffix _i
//               mod  C_1POINT0_ON  -> C_XCLIP_1POINT0
//151220su      :mk easy to inference ROM coding in MAX10
//              :mk easy to inference ROM coding in Cyclone I
//151218fr      : rm ~~~_inc.v
//                sin table +0.5
//                retruct external rom ~~~_inc.v
//151215tu      :mod selectanble to clip 1.0
//151213su      :1st.
module SIN_TBL_s11_s11 #(
        parameter C_XCLIP_1POINT0 = 0 //0: CLIP
                                      //1: non CLIP
)(
          CK_i
        , XARST_i
        , EN_CK_i
        , DAT_i   //2's -h800 0 +7FFF
        , SIN_o   //2's -h800 0 +h800
);

        localparam integer C_QQ_W = 
                (C_XCLIP_1POINT0 !=0) ? //0:clip 1:non clip
                        13
                :
                        12 
        ;

        input                           CK_i    ;
        input   tri0                    XARST_i ;
        input   tri1                    EN_CK_i ;
        input   tri0    [11 :0]         DAT_i     ; //2's -h800 0 +7FFF
        output          [C_QQ_W-1 :0]    SIN_o     ; //2's -h800 0 +h800
        // main
        wire    [ 9 :0] sin_adr         ;
        wire            down_curve      ;
        assign sin_adr = ( down_curve ) ? -DAT_i[ 9 :0] : DAT_i[9 :0] ;

        // 2CK_i dly
        wire    [ 8 :0] SIN_ROM_DAT     ;
        SIN_ROM_4s11_s11 u_SIN_ROM (
                  .CK_i         ( CK_i          )
                , .EN_CK_i      ( EN_CK_i       )
                , .ADR_i        ( sin_adr       )
                , .QQ_o         ( SIN_ROM_DAT   )
        ) ;
       
        reg     [ 9 :0] SIN_ADR_D     ;
        reg     [ 9 :0] SIN_ADR_DD    ;
        always @(posedge CK_i or negedge XARST_i) 
            if ( ~ XARST_i) begin
                SIN_ADR_D  <= 'd0 ;
                SIN_ADR_DD <= 'd0 ;
            end else if ( EN_CK_i) begin
                SIN_ADR_D  <= sin_adr ;
                SIN_ADR_DD <= SIN_ADR_D ;
            end
        wire    [12 :0] sin_dat ;
        assign sin_dat = SIN_ROM_DAT + {SIN_ADR_DD , 1'b0} ;

        reg             MINUS           ;
        reg             MAX_MIN         ;
        reg             ZERO            ;
        reg     [C_QQ_W-1 :0] SIN      ;
        always @ (posedge CK_i or negedge XARST_i)
                if ( ~ XARST_i ) begin
                        SIN <= 'd0 ;
                end else if (EN_CK_i) begin
                        if (C_XCLIP_1POINT0 != 0) begin //0:clip 1:non_clip
                                if ( ZERO )
                                        SIN <= 13'd0 ;
                                else if ( MAX_MIN )
                                        if ( MINUS )
                                                SIN <= -13'h800 ;
                                        else
                                                SIN <= 13'h800 ;
        
                                else
                                        if ( MINUS )
                                                SIN <= -sin_dat ;
                                        else
                                                SIN <= sin_dat ;
                        end else begin
                                if ( ZERO )
                                        SIN <= 12'd0 ;
                                else if (MAX_MIN | |sin_dat[12:11])
                                        if ( MINUS )
                                                SIN <= -12'h7FF ;
                                        else
                                                SIN <= 12'h7FF ;
                                else 
                                        if ( MINUS )
                                                SIN <= -sin_dat ;
                                        else
                                                SIN <= sin_dat ;
                        end
                end
        assign SIN_o = SIN ;


        // ctl
        assign down_curve = DAT_i[10] ;
        reg     MINUS_AD        ;
        reg     ZERO_AD         ;
        reg     MAX_MIN_AD      ;
        always @ (posedge CK_i or negedge XARST_i)
                if ( ~ XARST_i ) begin
                        MINUS_AD <= 1'b0 ;
                        MINUS <= 1'b0 ;
                        MAX_MIN_AD <= 1'b0 ;
                        MAX_MIN <= 1'b0 ;
                        ZERO_AD <= 1'b1 ;
                        ZERO <= 1'b1 ;
                end else if ( EN_CK_i) begin
                        MINUS_AD <= DAT_i[11] ;
                        MAX_MIN_AD <= (DAT_i[9:0] == 'd0) ;
                        ZERO_AD <= (DAT_i[9:0] == 'd0) & ~ DAT_i[10] ;
                        MINUS <= MINUS_AD ;
                        MAX_MIN <= MAX_MIN_AD ;
                        ZERO <= ZERO_AD ;
                end

endmodule // SIN_TBL_s11_s11

// 2ck dly
module SIN_ROM_4s11_s11 (
          CK_i
        , EN_CK_i
        , ADR_i
        , QQ_o
) ;
        input           CK_i      ;
        input           EN_CK_i ;
        input   [ 9 :0] ADR_i   ;
        output  [ 8 :0] QQ_o    ;


        reg     [ 9 :0] ROM_ADR ;
        always @ (posedge CK_i)
            if ( EN_CK_i )
                ROM_ADR <= ADR_i ;

//        `include "SIN_TBL_s11_s11_inc.v"
        // sin_tb_12_12_inc.v
        // datetime.datetime(2015, 12, 20, 11, 29, 28, 266222)
        reg    [ 8 :0] QQ     ;
        always @ (posedge CK_i)
            if ( EN_CK_i )
                case ( ROM_ADR )
                        10'h000 : QQ <= 9'h000 ;
                        10'h001 : QQ <= 9'h001 ;
                        10'h002 : QQ <= 9'h002 ;
                        10'h003 : QQ <= 9'h003 ;
                        10'h004 : QQ <= 9'h005 ;
                        10'h005 : QQ <= 9'h006 ;
                        10'h006 : QQ <= 9'h007 ;
                        10'h007 : QQ <= 9'h008 ;
                        10'h008 : QQ <= 9'h009 ;
                        10'h009 : QQ <= 9'h00A ;
                        10'h00A : QQ <= 9'h00B ;
                        10'h00B : QQ <= 9'h00D ;
                        10'h00C : QQ <= 9'h00E ;
                        10'h00D : QQ <= 9'h00F ;
                        10'h00E : QQ <= 9'h010 ;
                        10'h00F : QQ <= 9'h011 ;
                        10'h010 : QQ <= 9'h012 ;
                        10'h011 : QQ <= 9'h013 ;
                        10'h012 : QQ <= 9'h015 ;
                        10'h013 : QQ <= 9'h016 ;
                        10'h014 : QQ <= 9'h017 ;
                        10'h015 : QQ <= 9'h018 ;
                        10'h016 : QQ <= 9'h019 ;
                        10'h017 : QQ <= 9'h01A ;
                        10'h018 : QQ <= 9'h01B ;
                        10'h019 : QQ <= 9'h01D ;
                        10'h01A : QQ <= 9'h01E ;
                        10'h01B : QQ <= 9'h01F ;
                        10'h01C : QQ <= 9'h020 ;
                        10'h01D : QQ <= 9'h021 ;
                        10'h01E : QQ <= 9'h022 ;
                        10'h01F : QQ <= 9'h023 ;
                        10'h020 : QQ <= 9'h024 ;
                        10'h021 : QQ <= 9'h026 ;
                        10'h022 : QQ <= 9'h027 ;
                        10'h023 : QQ <= 9'h028 ;
                        10'h024 : QQ <= 9'h029 ;
                        10'h025 : QQ <= 9'h02A ;
                        10'h026 : QQ <= 9'h02B ;
                        10'h027 : QQ <= 9'h02C ;
                        10'h028 : QQ <= 9'h02E ;
                        10'h029 : QQ <= 9'h02F ;
                        10'h02A : QQ <= 9'h030 ;
                        10'h02B : QQ <= 9'h031 ;
                        10'h02C : QQ <= 9'h032 ;
                        10'h02D : QQ <= 9'h033 ;
                        10'h02E : QQ <= 9'h034 ;
                        10'h02F : QQ <= 9'h036 ;
                        10'h030 : QQ <= 9'h037 ;
                        10'h031 : QQ <= 9'h038 ;
                        10'h032 : QQ <= 9'h039 ;
                        10'h033 : QQ <= 9'h03A ;
                        10'h034 : QQ <= 9'h03B ;
                        10'h035 : QQ <= 9'h03C ;
                        10'h036 : QQ <= 9'h03D ;
                        10'h037 : QQ <= 9'h03F ;
                        10'h038 : QQ <= 9'h040 ;
                        10'h039 : QQ <= 9'h041 ;
                        10'h03A : QQ <= 9'h042 ;
                        10'h03B : QQ <= 9'h043 ;
                        10'h03C : QQ <= 9'h044 ;
                        10'h03D : QQ <= 9'h045 ;
                        10'h03E : QQ <= 9'h046 ;
                        10'h03F : QQ <= 9'h048 ;
                        10'h040 : QQ <= 9'h049 ;
                        10'h041 : QQ <= 9'h04A ;
                        10'h042 : QQ <= 9'h04B ;
                        10'h043 : QQ <= 9'h04C ;
                        10'h044 : QQ <= 9'h04D ;
                        10'h045 : QQ <= 9'h04E ;
                        10'h046 : QQ <= 9'h04F ;
                        10'h047 : QQ <= 9'h051 ;
                        10'h048 : QQ <= 9'h052 ;
                        10'h049 : QQ <= 9'h053 ;
                        10'h04A : QQ <= 9'h054 ;
                        10'h04B : QQ <= 9'h055 ;
                        10'h04C : QQ <= 9'h056 ;
                        10'h04D : QQ <= 9'h057 ;
                        10'h04E : QQ <= 9'h058 ;
                        10'h04F : QQ <= 9'h05A ;
                        10'h050 : QQ <= 9'h05B ;
                        10'h051 : QQ <= 9'h05C ;
                        10'h052 : QQ <= 9'h05D ;
                        10'h053 : QQ <= 9'h05E ;
                        10'h054 : QQ <= 9'h05F ;
                        10'h055 : QQ <= 9'h060 ;
                        10'h056 : QQ <= 9'h061 ;
                        10'h057 : QQ <= 9'h063 ;
                        10'h058 : QQ <= 9'h064 ;
                        10'h059 : QQ <= 9'h065 ;
                        10'h05A : QQ <= 9'h066 ;
                        10'h05B : QQ <= 9'h067 ;
                        10'h05C : QQ <= 9'h068 ;
                        10'h05D : QQ <= 9'h069 ;
                        10'h05E : QQ <= 9'h06A ;
                        10'h05F : QQ <= 9'h06B ;
                        10'h060 : QQ <= 9'h06D ;
                        10'h061 : QQ <= 9'h06E ;
                        10'h062 : QQ <= 9'h06F ;
                        10'h063 : QQ <= 9'h070 ;
                        10'h064 : QQ <= 9'h071 ;
                        10'h065 : QQ <= 9'h072 ;
                        10'h066 : QQ <= 9'h073 ;
                        10'h067 : QQ <= 9'h074 ;
                        10'h068 : QQ <= 9'h075 ;
                        10'h069 : QQ <= 9'h076 ;
                        10'h06A : QQ <= 9'h078 ;
                        10'h06B : QQ <= 9'h079 ;
                        10'h06C : QQ <= 9'h07A ;
                        10'h06D : QQ <= 9'h07B ;
                        10'h06E : QQ <= 9'h07C ;
                        10'h06F : QQ <= 9'h07D ;
                        10'h070 : QQ <= 9'h07E ;
                        10'h071 : QQ <= 9'h07F ;
                        10'h072 : QQ <= 9'h080 ;
                        10'h073 : QQ <= 9'h081 ;
                        10'h074 : QQ <= 9'h083 ;
                        10'h075 : QQ <= 9'h084 ;
                        10'h076 : QQ <= 9'h085 ;
                        10'h077 : QQ <= 9'h086 ;
                        10'h078 : QQ <= 9'h087 ;
                        10'h079 : QQ <= 9'h088 ;
                        10'h07A : QQ <= 9'h089 ;
                        10'h07B : QQ <= 9'h08A ;
                        10'h07C : QQ <= 9'h08B ;
                        10'h07D : QQ <= 9'h08C ;
                        10'h07E : QQ <= 9'h08D ;
                        10'h07F : QQ <= 9'h08E ;
                        10'h080 : QQ <= 9'h090 ;
                        10'h081 : QQ <= 9'h091 ;
                        10'h082 : QQ <= 9'h092 ;
                        10'h083 : QQ <= 9'h093 ;
                        10'h084 : QQ <= 9'h094 ;
                        10'h085 : QQ <= 9'h095 ;
                        10'h086 : QQ <= 9'h096 ;
                        10'h087 : QQ <= 9'h097 ;
                        10'h088 : QQ <= 9'h098 ;
                        10'h089 : QQ <= 9'h099 ;
                        10'h08A : QQ <= 9'h09A ;
                        10'h08B : QQ <= 9'h09B ;
                        10'h08C : QQ <= 9'h09C ;
                        10'h08D : QQ <= 9'h09E ;
                        10'h08E : QQ <= 9'h09F ;
                        10'h08F : QQ <= 9'h0A0 ;
                        10'h090 : QQ <= 9'h0A1 ;
                        10'h091 : QQ <= 9'h0A2 ;
                        10'h092 : QQ <= 9'h0A3 ;
                        10'h093 : QQ <= 9'h0A4 ;
                        10'h094 : QQ <= 9'h0A5 ;
                        10'h095 : QQ <= 9'h0A6 ;
                        10'h096 : QQ <= 9'h0A7 ;
                        10'h097 : QQ <= 9'h0A8 ;
                        10'h098 : QQ <= 9'h0A9 ;
                        10'h099 : QQ <= 9'h0AA ;
                        10'h09A : QQ <= 9'h0AB ;
                        10'h09B : QQ <= 9'h0AC ;
                        10'h09C : QQ <= 9'h0AD ;
                        10'h09D : QQ <= 9'h0AE ;
                        10'h09E : QQ <= 9'h0B0 ;
                        10'h09F : QQ <= 9'h0B1 ;
                        10'h0A0 : QQ <= 9'h0B2 ;
                        10'h0A1 : QQ <= 9'h0B3 ;
                        10'h0A2 : QQ <= 9'h0B4 ;
                        10'h0A3 : QQ <= 9'h0B5 ;
                        10'h0A4 : QQ <= 9'h0B6 ;
                        10'h0A5 : QQ <= 9'h0B7 ;
                        10'h0A6 : QQ <= 9'h0B8 ;
                        10'h0A7 : QQ <= 9'h0B9 ;
                        10'h0A8 : QQ <= 9'h0BA ;
                        10'h0A9 : QQ <= 9'h0BB ;
                        10'h0AA : QQ <= 9'h0BC ;
                        10'h0AB : QQ <= 9'h0BD ;
                        10'h0AC : QQ <= 9'h0BE ;
                        10'h0AD : QQ <= 9'h0BF ;
                        10'h0AE : QQ <= 9'h0C0 ;
                        10'h0AF : QQ <= 9'h0C1 ;
                        10'h0B0 : QQ <= 9'h0C2 ;
                        10'h0B1 : QQ <= 9'h0C3 ;
                        10'h0B2 : QQ <= 9'h0C4 ;
                        10'h0B3 : QQ <= 9'h0C5 ;
                        10'h0B4 : QQ <= 9'h0C6 ;
                        10'h0B5 : QQ <= 9'h0C7 ;
                        10'h0B6 : QQ <= 9'h0C8 ;
                        10'h0B7 : QQ <= 9'h0C9 ;
                        10'h0B8 : QQ <= 9'h0CA ;
                        10'h0B9 : QQ <= 9'h0CB ;
                        10'h0BA : QQ <= 9'h0CC ;
                        10'h0BB : QQ <= 9'h0CD ;
                        10'h0BC : QQ <= 9'h0CE ;
                        10'h0BD : QQ <= 9'h0CF ;
                        10'h0BE : QQ <= 9'h0D0 ;
                        10'h0BF : QQ <= 9'h0D1 ;
                        10'h0C0 : QQ <= 9'h0D3 ;
                        10'h0C1 : QQ <= 9'h0D4 ;
                        10'h0C2 : QQ <= 9'h0D5 ;
                        10'h0C3 : QQ <= 9'h0D6 ;
                        10'h0C4 : QQ <= 9'h0D7 ;
                        10'h0C5 : QQ <= 9'h0D8 ;
                        10'h0C6 : QQ <= 9'h0D9 ;
                        10'h0C7 : QQ <= 9'h0DA ;
                        10'h0C8 : QQ <= 9'h0DB ;
                        10'h0C9 : QQ <= 9'h0DC ;
                        10'h0CA : QQ <= 9'h0DC ;
                        10'h0CB : QQ <= 9'h0DD ;
                        10'h0CC : QQ <= 9'h0DE ;
                        10'h0CD : QQ <= 9'h0DF ;
                        10'h0CE : QQ <= 9'h0E0 ;
                        10'h0CF : QQ <= 9'h0E1 ;
                        10'h0D0 : QQ <= 9'h0E2 ;
                        10'h0D1 : QQ <= 9'h0E3 ;
                        10'h0D2 : QQ <= 9'h0E4 ;
                        10'h0D3 : QQ <= 9'h0E5 ;
                        10'h0D4 : QQ <= 9'h0E6 ;
                        10'h0D5 : QQ <= 9'h0E7 ;
                        10'h0D6 : QQ <= 9'h0E8 ;
                        10'h0D7 : QQ <= 9'h0E9 ;
                        10'h0D8 : QQ <= 9'h0EA ;
                        10'h0D9 : QQ <= 9'h0EB ;
                        10'h0DA : QQ <= 9'h0EC ;
                        10'h0DB : QQ <= 9'h0ED ;
                        10'h0DC : QQ <= 9'h0EE ;
                        10'h0DD : QQ <= 9'h0EF ;
                        10'h0DE : QQ <= 9'h0F0 ;
                        10'h0DF : QQ <= 9'h0F1 ;
                        10'h0E0 : QQ <= 9'h0F2 ;
                        10'h0E1 : QQ <= 9'h0F3 ;
                        10'h0E2 : QQ <= 9'h0F4 ;
                        10'h0E3 : QQ <= 9'h0F5 ;
                        10'h0E4 : QQ <= 9'h0F6 ;
                        10'h0E5 : QQ <= 9'h0F7 ;
                        10'h0E6 : QQ <= 9'h0F8 ;
                        10'h0E7 : QQ <= 9'h0F9 ;
                        10'h0E8 : QQ <= 9'h0FA ;
                        10'h0E9 : QQ <= 9'h0FB ;
                        10'h0EA : QQ <= 9'h0FB ;
                        10'h0EB : QQ <= 9'h0FC ;
                        10'h0EC : QQ <= 9'h0FD ;
                        10'h0ED : QQ <= 9'h0FE ;
                        10'h0EE : QQ <= 9'h0FF ;
                        10'h0EF : QQ <= 9'h100 ;
                        10'h0F0 : QQ <= 9'h101 ;
                        10'h0F1 : QQ <= 9'h102 ;
                        10'h0F2 : QQ <= 9'h103 ;
                        10'h0F3 : QQ <= 9'h104 ;
                        10'h0F4 : QQ <= 9'h105 ;
                        10'h0F5 : QQ <= 9'h106 ;
                        10'h0F6 : QQ <= 9'h107 ;
                        10'h0F7 : QQ <= 9'h108 ;
                        10'h0F8 : QQ <= 9'h108 ;
                        10'h0F9 : QQ <= 9'h109 ;
                        10'h0FA : QQ <= 9'h10A ;
                        10'h0FB : QQ <= 9'h10B ;
                        10'h0FC : QQ <= 9'h10C ;
                        10'h0FD : QQ <= 9'h10D ;
                        10'h0FE : QQ <= 9'h10E ;
                        10'h0FF : QQ <= 9'h10F ;
                        10'h100 : QQ <= 9'h110 ;
                        10'h101 : QQ <= 9'h111 ;
                        10'h102 : QQ <= 9'h112 ;
                        10'h103 : QQ <= 9'h112 ;
                        10'h104 : QQ <= 9'h113 ;
                        10'h105 : QQ <= 9'h114 ;
                        10'h106 : QQ <= 9'h115 ;
                        10'h107 : QQ <= 9'h116 ;
                        10'h108 : QQ <= 9'h117 ;
                        10'h109 : QQ <= 9'h118 ;
                        10'h10A : QQ <= 9'h119 ;
                        10'h10B : QQ <= 9'h11A ;
                        10'h10C : QQ <= 9'h11A ;
                        10'h10D : QQ <= 9'h11B ;
                        10'h10E : QQ <= 9'h11C ;
                        10'h10F : QQ <= 9'h11D ;
                        10'h110 : QQ <= 9'h11E ;
                        10'h111 : QQ <= 9'h11F ;
                        10'h112 : QQ <= 9'h120 ;
                        10'h113 : QQ <= 9'h121 ;
                        10'h114 : QQ <= 9'h121 ;
                        10'h115 : QQ <= 9'h122 ;
                        10'h116 : QQ <= 9'h123 ;
                        10'h117 : QQ <= 9'h124 ;
                        10'h118 : QQ <= 9'h125 ;
                        10'h119 : QQ <= 9'h126 ;
                        10'h11A : QQ <= 9'h127 ;
                        10'h11B : QQ <= 9'h127 ;
                        10'h11C : QQ <= 9'h128 ;
                        10'h11D : QQ <= 9'h129 ;
                        10'h11E : QQ <= 9'h12A ;
                        10'h11F : QQ <= 9'h12B ;
                        10'h120 : QQ <= 9'h12C ;
                        10'h121 : QQ <= 9'h12C ;
                        10'h122 : QQ <= 9'h12D ;
                        10'h123 : QQ <= 9'h12E ;
                        10'h124 : QQ <= 9'h12F ;
                        10'h125 : QQ <= 9'h130 ;
                        10'h126 : QQ <= 9'h131 ;
                        10'h127 : QQ <= 9'h131 ;
                        10'h128 : QQ <= 9'h132 ;
                        10'h129 : QQ <= 9'h133 ;
                        10'h12A : QQ <= 9'h134 ;
                        10'h12B : QQ <= 9'h135 ;
                        10'h12C : QQ <= 9'h136 ;
                        10'h12D : QQ <= 9'h136 ;
                        10'h12E : QQ <= 9'h137 ;
                        10'h12F : QQ <= 9'h138 ;
                        10'h130 : QQ <= 9'h139 ;
                        10'h131 : QQ <= 9'h13A ;
                        10'h132 : QQ <= 9'h13A ;
                        10'h133 : QQ <= 9'h13B ;
                        10'h134 : QQ <= 9'h13C ;
                        10'h135 : QQ <= 9'h13D ;
                        10'h136 : QQ <= 9'h13E ;
                        10'h137 : QQ <= 9'h13E ;
                        10'h138 : QQ <= 9'h13F ;
                        10'h139 : QQ <= 9'h140 ;
                        10'h13A : QQ <= 9'h141 ;
                        10'h13B : QQ <= 9'h142 ;
                        10'h13C : QQ <= 9'h142 ;
                        10'h13D : QQ <= 9'h143 ;
                        10'h13E : QQ <= 9'h144 ;
                        10'h13F : QQ <= 9'h145 ;
                        10'h140 : QQ <= 9'h145 ;
                        10'h141 : QQ <= 9'h146 ;
                        10'h142 : QQ <= 9'h147 ;
                        10'h143 : QQ <= 9'h148 ;
                        10'h144 : QQ <= 9'h148 ;
                        10'h145 : QQ <= 9'h149 ;
                        10'h146 : QQ <= 9'h14A ;
                        10'h147 : QQ <= 9'h14B ;
                        10'h148 : QQ <= 9'h14C ;
                        10'h149 : QQ <= 9'h14C ;
                        10'h14A : QQ <= 9'h14D ;
                        10'h14B : QQ <= 9'h14E ;
                        10'h14C : QQ <= 9'h14F ;
                        10'h14D : QQ <= 9'h14F ;
                        10'h14E : QQ <= 9'h150 ;
                        10'h14F : QQ <= 9'h151 ;
                        10'h150 : QQ <= 9'h151 ;
                        10'h151 : QQ <= 9'h152 ;
                        10'h152 : QQ <= 9'h153 ;
                        10'h153 : QQ <= 9'h154 ;
                        10'h154 : QQ <= 9'h154 ;
                        10'h155 : QQ <= 9'h155 ;
                        10'h156 : QQ <= 9'h156 ;
                        10'h157 : QQ <= 9'h157 ;
                        10'h158 : QQ <= 9'h157 ;
                        10'h159 : QQ <= 9'h158 ;
                        10'h15A : QQ <= 9'h159 ;
                        10'h15B : QQ <= 9'h159 ;
                        10'h15C : QQ <= 9'h15A ;
                        10'h15D : QQ <= 9'h15B ;
                        10'h15E : QQ <= 9'h15B ;
                        10'h15F : QQ <= 9'h15C ;
                        10'h160 : QQ <= 9'h15D ;
                        10'h161 : QQ <= 9'h15E ;
                        10'h162 : QQ <= 9'h15E ;
                        10'h163 : QQ <= 9'h15F ;
                        10'h164 : QQ <= 9'h160 ;
                        10'h165 : QQ <= 9'h160 ;
                        10'h166 : QQ <= 9'h161 ;
                        10'h167 : QQ <= 9'h162 ;
                        10'h168 : QQ <= 9'h162 ;
                        10'h169 : QQ <= 9'h163 ;
                        10'h16A : QQ <= 9'h164 ;
                        10'h16B : QQ <= 9'h164 ;
                        10'h16C : QQ <= 9'h165 ;
                        10'h16D : QQ <= 9'h166 ;
                        10'h16E : QQ <= 9'h166 ;
                        10'h16F : QQ <= 9'h167 ;
                        10'h170 : QQ <= 9'h168 ;
                        10'h171 : QQ <= 9'h168 ;
                        10'h172 : QQ <= 9'h169 ;
                        10'h173 : QQ <= 9'h16A ;
                        10'h174 : QQ <= 9'h16A ;
                        10'h175 : QQ <= 9'h16B ;
                        10'h176 : QQ <= 9'h16C ;
                        10'h177 : QQ <= 9'h16C ;
                        10'h178 : QQ <= 9'h16D ;
                        10'h179 : QQ <= 9'h16D ;
                        10'h17A : QQ <= 9'h16E ;
                        10'h17B : QQ <= 9'h16F ;
                        10'h17C : QQ <= 9'h16F ;
                        10'h17D : QQ <= 9'h170 ;
                        10'h17E : QQ <= 9'h171 ;
                        10'h17F : QQ <= 9'h171 ;
                        10'h180 : QQ <= 9'h172 ;
                        10'h181 : QQ <= 9'h172 ;
                        10'h182 : QQ <= 9'h173 ;
                        10'h183 : QQ <= 9'h174 ;
                        10'h184 : QQ <= 9'h174 ;
                        10'h185 : QQ <= 9'h175 ;
                        10'h186 : QQ <= 9'h175 ;
                        10'h187 : QQ <= 9'h176 ;
                        10'h188 : QQ <= 9'h177 ;
                        10'h189 : QQ <= 9'h177 ;
                        10'h18A : QQ <= 9'h178 ;
                        10'h18B : QQ <= 9'h178 ;
                        10'h18C : QQ <= 9'h179 ;
                        10'h18D : QQ <= 9'h17A ;
                        10'h18E : QQ <= 9'h17A ;
                        10'h18F : QQ <= 9'h17B ;
                        10'h190 : QQ <= 9'h17B ;
                        10'h191 : QQ <= 9'h17C ;
                        10'h192 : QQ <= 9'h17C ;
                        10'h193 : QQ <= 9'h17D ;
                        10'h194 : QQ <= 9'h17E ;
                        10'h195 : QQ <= 9'h17E ;
                        10'h196 : QQ <= 9'h17F ;
                        10'h197 : QQ <= 9'h17F ;
                        10'h198 : QQ <= 9'h180 ;
                        10'h199 : QQ <= 9'h180 ;
                        10'h19A : QQ <= 9'h181 ;
                        10'h19B : QQ <= 9'h181 ;
                        10'h19C : QQ <= 9'h182 ;
                        10'h19D : QQ <= 9'h182 ;
                        10'h19E : QQ <= 9'h183 ;
                        10'h19F : QQ <= 9'h183 ;
                        10'h1A0 : QQ <= 9'h184 ;
                        10'h1A1 : QQ <= 9'h185 ;
                        10'h1A2 : QQ <= 9'h185 ;
                        10'h1A3 : QQ <= 9'h186 ;
                        10'h1A4 : QQ <= 9'h186 ;
                        10'h1A5 : QQ <= 9'h187 ;
                        10'h1A6 : QQ <= 9'h187 ;
                        10'h1A7 : QQ <= 9'h188 ;
                        10'h1A8 : QQ <= 9'h188 ;
                        10'h1A9 : QQ <= 9'h189 ;
                        10'h1AA : QQ <= 9'h189 ;
                        10'h1AB : QQ <= 9'h18A ;
                        10'h1AC : QQ <= 9'h18A ;
                        10'h1AD : QQ <= 9'h18B ;
                        10'h1AE : QQ <= 9'h18B ;
                        10'h1AF : QQ <= 9'h18C ;
                        10'h1B0 : QQ <= 9'h18C ;
                        10'h1B1 : QQ <= 9'h18C ;
                        10'h1B2 : QQ <= 9'h18D ;
                        10'h1B3 : QQ <= 9'h18D ;
                        10'h1B4 : QQ <= 9'h18E ;
                        10'h1B5 : QQ <= 9'h18E ;
                        10'h1B6 : QQ <= 9'h18F ;
                        10'h1B7 : QQ <= 9'h18F ;
                        10'h1B8 : QQ <= 9'h190 ;
                        10'h1B9 : QQ <= 9'h190 ;
                        10'h1BA : QQ <= 9'h191 ;
                        10'h1BB : QQ <= 9'h191 ;
                        10'h1BC : QQ <= 9'h191 ;
                        10'h1BD : QQ <= 9'h192 ;
                        10'h1BE : QQ <= 9'h192 ;
                        10'h1BF : QQ <= 9'h193 ;
                        10'h1C0 : QQ <= 9'h193 ;
                        10'h1C1 : QQ <= 9'h194 ;
                        10'h1C2 : QQ <= 9'h194 ;
                        10'h1C3 : QQ <= 9'h195 ;
                        10'h1C4 : QQ <= 9'h195 ;
                        10'h1C5 : QQ <= 9'h195 ;
                        10'h1C6 : QQ <= 9'h196 ;
                        10'h1C7 : QQ <= 9'h196 ;
                        10'h1C8 : QQ <= 9'h197 ;
                        10'h1C9 : QQ <= 9'h197 ;
                        10'h1CA : QQ <= 9'h197 ;
                        10'h1CB : QQ <= 9'h198 ;
                        10'h1CC : QQ <= 9'h198 ;
                        10'h1CD : QQ <= 9'h199 ;
                        10'h1CE : QQ <= 9'h199 ;
                        10'h1CF : QQ <= 9'h199 ;
                        10'h1D0 : QQ <= 9'h19A ;
                        10'h1D1 : QQ <= 9'h19A ;
                        10'h1D2 : QQ <= 9'h19A ;
                        10'h1D3 : QQ <= 9'h19B ;
                        10'h1D4 : QQ <= 9'h19B ;
                        10'h1D5 : QQ <= 9'h19C ;
                        10'h1D6 : QQ <= 9'h19C ;
                        10'h1D7 : QQ <= 9'h19C ;
                        10'h1D8 : QQ <= 9'h19D ;
                        10'h1D9 : QQ <= 9'h19D ;
                        10'h1DA : QQ <= 9'h19D ;
                        10'h1DB : QQ <= 9'h19E ;
                        10'h1DC : QQ <= 9'h19E ;
                        10'h1DD : QQ <= 9'h19E ;
                        10'h1DE : QQ <= 9'h19F ;
                        10'h1DF : QQ <= 9'h19F ;
                        10'h1E0 : QQ <= 9'h19F ;
                        10'h1E1 : QQ <= 9'h1A0 ;
                        10'h1E2 : QQ <= 9'h1A0 ;
                        10'h1E3 : QQ <= 9'h1A0 ;
                        10'h1E4 : QQ <= 9'h1A1 ;
                        10'h1E5 : QQ <= 9'h1A1 ;
                        10'h1E6 : QQ <= 9'h1A1 ;
                        10'h1E7 : QQ <= 9'h1A2 ;
                        10'h1E8 : QQ <= 9'h1A2 ;
                        10'h1E9 : QQ <= 9'h1A2 ;
                        10'h1EA : QQ <= 9'h1A2 ;
                        10'h1EB : QQ <= 9'h1A3 ;
                        10'h1EC : QQ <= 9'h1A3 ;
                        10'h1ED : QQ <= 9'h1A3 ;
                        10'h1EE : QQ <= 9'h1A4 ;
                        10'h1EF : QQ <= 9'h1A4 ;
                        10'h1F0 : QQ <= 9'h1A4 ;
                        10'h1F1 : QQ <= 9'h1A4 ;
                        10'h1F2 : QQ <= 9'h1A5 ;
                        10'h1F3 : QQ <= 9'h1A5 ;
                        10'h1F4 : QQ <= 9'h1A5 ;
                        10'h1F5 : QQ <= 9'h1A6 ;
                        10'h1F6 : QQ <= 9'h1A6 ;
                        10'h1F7 : QQ <= 9'h1A6 ;
                        10'h1F8 : QQ <= 9'h1A6 ;
                        10'h1F9 : QQ <= 9'h1A7 ;
                        10'h1FA : QQ <= 9'h1A7 ;
                        10'h1FB : QQ <= 9'h1A7 ;
                        10'h1FC : QQ <= 9'h1A7 ;
                        10'h1FD : QQ <= 9'h1A7 ;
                        10'h1FE : QQ <= 9'h1A8 ;
                        10'h1FF : QQ <= 9'h1A8 ;
                        10'h200 : QQ <= 9'h1A8 ;
                        10'h201 : QQ <= 9'h1A8 ;
                        10'h202 : QQ <= 9'h1A9 ;
                        10'h203 : QQ <= 9'h1A9 ;
                        10'h204 : QQ <= 9'h1A9 ;
                        10'h205 : QQ <= 9'h1A9 ;
                        10'h206 : QQ <= 9'h1A9 ;
                        10'h207 : QQ <= 9'h1AA ;
                        10'h208 : QQ <= 9'h1AA ;
                        10'h209 : QQ <= 9'h1AA ;
                        10'h20A : QQ <= 9'h1AA ;
                        10'h20B : QQ <= 9'h1AA ;
                        10'h20C : QQ <= 9'h1AB ;
                        10'h20D : QQ <= 9'h1AB ;
                        10'h20E : QQ <= 9'h1AB ;
                        10'h20F : QQ <= 9'h1AB ;
                        10'h210 : QQ <= 9'h1AB ;
                        10'h211 : QQ <= 9'h1AB ;
                        10'h212 : QQ <= 9'h1AC ;
                        10'h213 : QQ <= 9'h1AC ;
                        10'h214 : QQ <= 9'h1AC ;
                        10'h215 : QQ <= 9'h1AC ;
                        10'h216 : QQ <= 9'h1AC ;
                        10'h217 : QQ <= 9'h1AC ;
                        10'h218 : QQ <= 9'h1AC ;
                        10'h219 : QQ <= 9'h1AD ;
                        10'h21A : QQ <= 9'h1AD ;
                        10'h21B : QQ <= 9'h1AD ;
                        10'h21C : QQ <= 9'h1AD ;
                        10'h21D : QQ <= 9'h1AD ;
                        10'h21E : QQ <= 9'h1AD ;
                        10'h21F : QQ <= 9'h1AD ;
                        10'h220 : QQ <= 9'h1AD ;
                        10'h221 : QQ <= 9'h1AE ;
                        10'h222 : QQ <= 9'h1AE ;
                        10'h223 : QQ <= 9'h1AE ;
                        10'h224 : QQ <= 9'h1AE ;
                        10'h225 : QQ <= 9'h1AE ;
                        10'h226 : QQ <= 9'h1AE ;
                        10'h227 : QQ <= 9'h1AE ;
                        10'h228 : QQ <= 9'h1AE ;
                        10'h229 : QQ <= 9'h1AE ;
                        10'h22A : QQ <= 9'h1AE ;
                        10'h22B : QQ <= 9'h1AE ;
                        10'h22C : QQ <= 9'h1AF ;
                        10'h22D : QQ <= 9'h1AF ;
                        10'h22E : QQ <= 9'h1AF ;
                        10'h22F : QQ <= 9'h1AF ;
                        10'h230 : QQ <= 9'h1AF ;
                        10'h231 : QQ <= 9'h1AF ;
                        10'h232 : QQ <= 9'h1AF ;
                        10'h233 : QQ <= 9'h1AF ;
                        10'h234 : QQ <= 9'h1AF ;
                        10'h235 : QQ <= 9'h1AF ;
                        10'h236 : QQ <= 9'h1AF ;
                        10'h237 : QQ <= 9'h1AF ;
                        10'h238 : QQ <= 9'h1AF ;
                        10'h239 : QQ <= 9'h1AF ;
                        10'h23A : QQ <= 9'h1AF ;
                        10'h23B : QQ <= 9'h1AF ;
                        10'h23C : QQ <= 9'h1AF ;
                        10'h23D : QQ <= 9'h1AF ;
                        10'h23E : QQ <= 9'h1AF ;
                        10'h23F : QQ <= 9'h1AF ;
                        10'h240 : QQ <= 9'h1AF ;
                        10'h241 : QQ <= 9'h1AF ;
                        10'h242 : QQ <= 9'h1AF ;
                        10'h243 : QQ <= 9'h1AF ;
                        10'h244 : QQ <= 9'h1AF ;
                        10'h245 : QQ <= 9'h1AF ;
                        10'h246 : QQ <= 9'h1AF ;
                        10'h247 : QQ <= 9'h1AF ;
                        10'h248 : QQ <= 9'h1AF ;
                        10'h249 : QQ <= 9'h1AF ;
                        10'h24A : QQ <= 9'h1AF ;
                        10'h24B : QQ <= 9'h1AF ;
                        10'h24C : QQ <= 9'h1AF ;
                        10'h24D : QQ <= 9'h1AF ;
                        10'h24E : QQ <= 9'h1AF ;
                        10'h24F : QQ <= 9'h1AF ;
                        10'h250 : QQ <= 9'h1AF ;
                        10'h251 : QQ <= 9'h1AE ;
                        10'h252 : QQ <= 9'h1AE ;
                        10'h253 : QQ <= 9'h1AE ;
                        10'h254 : QQ <= 9'h1AE ;
                        10'h255 : QQ <= 9'h1AE ;
                        10'h256 : QQ <= 9'h1AE ;
                        10'h257 : QQ <= 9'h1AE ;
                        10'h258 : QQ <= 9'h1AE ;
                        10'h259 : QQ <= 9'h1AE ;
                        10'h25A : QQ <= 9'h1AE ;
                        10'h25B : QQ <= 9'h1AE ;
                        10'h25C : QQ <= 9'h1AD ;
                        10'h25D : QQ <= 9'h1AD ;
                        10'h25E : QQ <= 9'h1AD ;
                        10'h25F : QQ <= 9'h1AD ;
                        10'h260 : QQ <= 9'h1AD ;
                        10'h261 : QQ <= 9'h1AD ;
                        10'h262 : QQ <= 9'h1AD ;
                        10'h263 : QQ <= 9'h1AD ;
                        10'h264 : QQ <= 9'h1AC ;
                        10'h265 : QQ <= 9'h1AC ;
                        10'h266 : QQ <= 9'h1AC ;
                        10'h267 : QQ <= 9'h1AC ;
                        10'h268 : QQ <= 9'h1AC ;
                        10'h269 : QQ <= 9'h1AC ;
                        10'h26A : QQ <= 9'h1AB ;
                        10'h26B : QQ <= 9'h1AB ;
                        10'h26C : QQ <= 9'h1AB ;
                        10'h26D : QQ <= 9'h1AB ;
                        10'h26E : QQ <= 9'h1AB ;
                        10'h26F : QQ <= 9'h1AB ;
                        10'h270 : QQ <= 9'h1AA ;
                        10'h271 : QQ <= 9'h1AA ;
                        10'h272 : QQ <= 9'h1AA ;
                        10'h273 : QQ <= 9'h1AA ;
                        10'h274 : QQ <= 9'h1AA ;
                        10'h275 : QQ <= 9'h1A9 ;
                        10'h276 : QQ <= 9'h1A9 ;
                        10'h277 : QQ <= 9'h1A9 ;
                        10'h278 : QQ <= 9'h1A9 ;
                        10'h279 : QQ <= 9'h1A9 ;
                        10'h27A : QQ <= 9'h1A8 ;
                        10'h27B : QQ <= 9'h1A8 ;
                        10'h27C : QQ <= 9'h1A8 ;
                        10'h27D : QQ <= 9'h1A8 ;
                        10'h27E : QQ <= 9'h1A7 ;
                        10'h27F : QQ <= 9'h1A7 ;
                        10'h280 : QQ <= 9'h1A7 ;
                        10'h281 : QQ <= 9'h1A7 ;
                        10'h282 : QQ <= 9'h1A6 ;
                        10'h283 : QQ <= 9'h1A6 ;
                        10'h284 : QQ <= 9'h1A6 ;
                        10'h285 : QQ <= 9'h1A6 ;
                        10'h286 : QQ <= 9'h1A5 ;
                        10'h287 : QQ <= 9'h1A5 ;
                        10'h288 : QQ <= 9'h1A5 ;
                        10'h289 : QQ <= 9'h1A4 ;
                        10'h28A : QQ <= 9'h1A4 ;
                        10'h28B : QQ <= 9'h1A4 ;
                        10'h28C : QQ <= 9'h1A4 ;
                        10'h28D : QQ <= 9'h1A3 ;
                        10'h28E : QQ <= 9'h1A3 ;
                        10'h28F : QQ <= 9'h1A3 ;
                        10'h290 : QQ <= 9'h1A2 ;
                        10'h291 : QQ <= 9'h1A2 ;
                        10'h292 : QQ <= 9'h1A2 ;
                        10'h293 : QQ <= 9'h1A1 ;
                        10'h294 : QQ <= 9'h1A1 ;
                        10'h295 : QQ <= 9'h1A1 ;
                        10'h296 : QQ <= 9'h1A0 ;
                        10'h297 : QQ <= 9'h1A0 ;
                        10'h298 : QQ <= 9'h1A0 ;
                        10'h299 : QQ <= 9'h19F ;
                        10'h29A : QQ <= 9'h19F ;
                        10'h29B : QQ <= 9'h19F ;
                        10'h29C : QQ <= 9'h19E ;
                        10'h29D : QQ <= 9'h19E ;
                        10'h29E : QQ <= 9'h19D ;
                        10'h29F : QQ <= 9'h19D ;
                        10'h2A0 : QQ <= 9'h19D ;
                        10'h2A1 : QQ <= 9'h19C ;
                        10'h2A2 : QQ <= 9'h19C ;
                        10'h2A3 : QQ <= 9'h19B ;
                        10'h2A4 : QQ <= 9'h19B ;
                        10'h2A5 : QQ <= 9'h19B ;
                        10'h2A6 : QQ <= 9'h19A ;
                        10'h2A7 : QQ <= 9'h19A ;
                        10'h2A8 : QQ <= 9'h199 ;
                        10'h2A9 : QQ <= 9'h199 ;
                        10'h2AA : QQ <= 9'h199 ;
                        10'h2AB : QQ <= 9'h198 ;
                        10'h2AC : QQ <= 9'h198 ;
                        10'h2AD : QQ <= 9'h197 ;
                        10'h2AE : QQ <= 9'h197 ;
                        10'h2AF : QQ <= 9'h196 ;
                        10'h2B0 : QQ <= 9'h196 ;
                        10'h2B1 : QQ <= 9'h195 ;
                        10'h2B2 : QQ <= 9'h195 ;
                        10'h2B3 : QQ <= 9'h195 ;
                        10'h2B4 : QQ <= 9'h194 ;
                        10'h2B5 : QQ <= 9'h194 ;
                        10'h2B6 : QQ <= 9'h193 ;
                        10'h2B7 : QQ <= 9'h193 ;
                        10'h2B8 : QQ <= 9'h192 ;
                        10'h2B9 : QQ <= 9'h192 ;
                        10'h2BA : QQ <= 9'h191 ;
                        10'h2BB : QQ <= 9'h191 ;
                        10'h2BC : QQ <= 9'h190 ;
                        10'h2BD : QQ <= 9'h190 ;
                        10'h2BE : QQ <= 9'h18F ;
                        10'h2BF : QQ <= 9'h18F ;
                        10'h2C0 : QQ <= 9'h18E ;
                        10'h2C1 : QQ <= 9'h18E ;
                        10'h2C2 : QQ <= 9'h18D ;
                        10'h2C3 : QQ <= 9'h18D ;
                        10'h2C4 : QQ <= 9'h18C ;
                        10'h2C5 : QQ <= 9'h18C ;
                        10'h2C6 : QQ <= 9'h18B ;
                        10'h2C7 : QQ <= 9'h18A ;
                        10'h2C8 : QQ <= 9'h18A ;
                        10'h2C9 : QQ <= 9'h189 ;
                        10'h2CA : QQ <= 9'h189 ;
                        10'h2CB : QQ <= 9'h188 ;
                        10'h2CC : QQ <= 9'h188 ;
                        10'h2CD : QQ <= 9'h187 ;
                        10'h2CE : QQ <= 9'h186 ;
                        10'h2CF : QQ <= 9'h186 ;
                        10'h2D0 : QQ <= 9'h185 ;
                        10'h2D1 : QQ <= 9'h185 ;
                        10'h2D2 : QQ <= 9'h184 ;
                        10'h2D3 : QQ <= 9'h184 ;
                        10'h2D4 : QQ <= 9'h183 ;
                        10'h2D5 : QQ <= 9'h182 ;
                        10'h2D6 : QQ <= 9'h182 ;
                        10'h2D7 : QQ <= 9'h181 ;
                        10'h2D8 : QQ <= 9'h180 ;
                        10'h2D9 : QQ <= 9'h180 ;
                        10'h2DA : QQ <= 9'h17F ;
                        10'h2DB : QQ <= 9'h17F ;
                        10'h2DC : QQ <= 9'h17E ;
                        10'h2DD : QQ <= 9'h17D ;
                        10'h2DE : QQ <= 9'h17D ;
                        10'h2DF : QQ <= 9'h17C ;
                        10'h2E0 : QQ <= 9'h17B ;
                        10'h2E1 : QQ <= 9'h17B ;
                        10'h2E2 : QQ <= 9'h17A ;
                        10'h2E3 : QQ <= 9'h179 ;
                        10'h2E4 : QQ <= 9'h179 ;
                        10'h2E5 : QQ <= 9'h178 ;
                        10'h2E6 : QQ <= 9'h177 ;
                        10'h2E7 : QQ <= 9'h177 ;
                        10'h2E8 : QQ <= 9'h176 ;
                        10'h2E9 : QQ <= 9'h175 ;
                        10'h2EA : QQ <= 9'h175 ;
                        10'h2EB : QQ <= 9'h174 ;
                        10'h2EC : QQ <= 9'h173 ;
                        10'h2ED : QQ <= 9'h172 ;
                        10'h2EE : QQ <= 9'h172 ;
                        10'h2EF : QQ <= 9'h171 ;
                        10'h2F0 : QQ <= 9'h170 ;
                        10'h2F1 : QQ <= 9'h170 ;
                        10'h2F2 : QQ <= 9'h16F ;
                        10'h2F3 : QQ <= 9'h16E ;
                        10'h2F4 : QQ <= 9'h16D ;
                        10'h2F5 : QQ <= 9'h16D ;
                        10'h2F6 : QQ <= 9'h16C ;
                        10'h2F7 : QQ <= 9'h16B ;
                        10'h2F8 : QQ <= 9'h16A ;
                        10'h2F9 : QQ <= 9'h16A ;
                        10'h2FA : QQ <= 9'h169 ;
                        10'h2FB : QQ <= 9'h168 ;
                        10'h2FC : QQ <= 9'h167 ;
                        10'h2FD : QQ <= 9'h166 ;
                        10'h2FE : QQ <= 9'h166 ;
                        10'h2FF : QQ <= 9'h165 ;
                        10'h300 : QQ <= 9'h164 ;
                        10'h301 : QQ <= 9'h163 ;
                        10'h302 : QQ <= 9'h163 ;
                        10'h303 : QQ <= 9'h162 ;
                        10'h304 : QQ <= 9'h161 ;
                        10'h305 : QQ <= 9'h160 ;
                        10'h306 : QQ <= 9'h15F ;
                        10'h307 : QQ <= 9'h15E ;
                        10'h308 : QQ <= 9'h15E ;
                        10'h309 : QQ <= 9'h15D ;
                        10'h30A : QQ <= 9'h15C ;
                        10'h30B : QQ <= 9'h15B ;
                        10'h30C : QQ <= 9'h15A ;
                        10'h30D : QQ <= 9'h159 ;
                        10'h30E : QQ <= 9'h158 ;
                        10'h30F : QQ <= 9'h158 ;
                        10'h310 : QQ <= 9'h157 ;
                        10'h311 : QQ <= 9'h156 ;
                        10'h312 : QQ <= 9'h155 ;
                        10'h313 : QQ <= 9'h154 ;
                        10'h314 : QQ <= 9'h153 ;
                        10'h315 : QQ <= 9'h152 ;
                        10'h316 : QQ <= 9'h151 ;
                        10'h317 : QQ <= 9'h151 ;
                        10'h318 : QQ <= 9'h150 ;
                        10'h319 : QQ <= 9'h14F ;
                        10'h31A : QQ <= 9'h14E ;
                        10'h31B : QQ <= 9'h14D ;
                        10'h31C : QQ <= 9'h14C ;
                        10'h31D : QQ <= 9'h14B ;
                        10'h31E : QQ <= 9'h14A ;
                        10'h31F : QQ <= 9'h149 ;
                        10'h320 : QQ <= 9'h148 ;
                        10'h321 : QQ <= 9'h147 ;
                        10'h322 : QQ <= 9'h146 ;
                        10'h323 : QQ <= 9'h145 ;
                        10'h324 : QQ <= 9'h144 ;
                        10'h325 : QQ <= 9'h144 ;
                        10'h326 : QQ <= 9'h143 ;
                        10'h327 : QQ <= 9'h142 ;
                        10'h328 : QQ <= 9'h141 ;
                        10'h329 : QQ <= 9'h140 ;
                        10'h32A : QQ <= 9'h13F ;
                        10'h32B : QQ <= 9'h13E ;
                        10'h32C : QQ <= 9'h13D ;
                        10'h32D : QQ <= 9'h13C ;
                        10'h32E : QQ <= 9'h13B ;
                        10'h32F : QQ <= 9'h13A ;
                        10'h330 : QQ <= 9'h139 ;
                        10'h331 : QQ <= 9'h138 ;
                        10'h332 : QQ <= 9'h137 ;
                        10'h333 : QQ <= 9'h136 ;
                        10'h334 : QQ <= 9'h135 ;
                        10'h335 : QQ <= 9'h134 ;
                        10'h336 : QQ <= 9'h132 ;
                        10'h337 : QQ <= 9'h131 ;
                        10'h338 : QQ <= 9'h130 ;
                        10'h339 : QQ <= 9'h12F ;
                        10'h33A : QQ <= 9'h12E ;
                        10'h33B : QQ <= 9'h12D ;
                        10'h33C : QQ <= 9'h12C ;
                        10'h33D : QQ <= 9'h12B ;
                        10'h33E : QQ <= 9'h12A ;
                        10'h33F : QQ <= 9'h129 ;
                        10'h340 : QQ <= 9'h128 ;
                        10'h341 : QQ <= 9'h127 ;
                        10'h342 : QQ <= 9'h126 ;
                        10'h343 : QQ <= 9'h125 ;
                        10'h344 : QQ <= 9'h123 ;
                        10'h345 : QQ <= 9'h122 ;
                        10'h346 : QQ <= 9'h121 ;
                        10'h347 : QQ <= 9'h120 ;
                        10'h348 : QQ <= 9'h11F ;
                        10'h349 : QQ <= 9'h11E ;
                        10'h34A : QQ <= 9'h11D ;
                        10'h34B : QQ <= 9'h11C ;
                        10'h34C : QQ <= 9'h11A ;
                        10'h34D : QQ <= 9'h119 ;
                        10'h34E : QQ <= 9'h118 ;
                        10'h34F : QQ <= 9'h117 ;
                        10'h350 : QQ <= 9'h116 ;
                        10'h351 : QQ <= 9'h115 ;
                        10'h352 : QQ <= 9'h113 ;
                        10'h353 : QQ <= 9'h112 ;
                        10'h354 : QQ <= 9'h111 ;
                        10'h355 : QQ <= 9'h110 ;
                        10'h356 : QQ <= 9'h10F ;
                        10'h357 : QQ <= 9'h10E ;
                        10'h358 : QQ <= 9'h10C ;
                        10'h359 : QQ <= 9'h10B ;
                        10'h35A : QQ <= 9'h10A ;
                        10'h35B : QQ <= 9'h109 ;
                        10'h35C : QQ <= 9'h108 ;
                        10'h35D : QQ <= 9'h106 ;
                        10'h35E : QQ <= 9'h105 ;
                        10'h35F : QQ <= 9'h104 ;
                        10'h360 : QQ <= 9'h103 ;
                        10'h361 : QQ <= 9'h101 ;
                        10'h362 : QQ <= 9'h100 ;
                        10'h363 : QQ <= 9'h0FF ;
                        10'h364 : QQ <= 9'h0FE ;
                        10'h365 : QQ <= 9'h0FC ;
                        10'h366 : QQ <= 9'h0FB ;
                        10'h367 : QQ <= 9'h0FA ;
                        10'h368 : QQ <= 9'h0F9 ;
                        10'h369 : QQ <= 9'h0F7 ;
                        10'h36A : QQ <= 9'h0F6 ;
                        10'h36B : QQ <= 9'h0F5 ;
                        10'h36C : QQ <= 9'h0F3 ;
                        10'h36D : QQ <= 9'h0F2 ;
                        10'h36E : QQ <= 9'h0F1 ;
                        10'h36F : QQ <= 9'h0F0 ;
                        10'h370 : QQ <= 9'h0EE ;
                        10'h371 : QQ <= 9'h0ED ;
                        10'h372 : QQ <= 9'h0EC ;
                        10'h373 : QQ <= 9'h0EA ;
                        10'h374 : QQ <= 9'h0E9 ;
                        10'h375 : QQ <= 9'h0E8 ;
                        10'h376 : QQ <= 9'h0E6 ;
                        10'h377 : QQ <= 9'h0E5 ;
                        10'h378 : QQ <= 9'h0E4 ;
                        10'h379 : QQ <= 9'h0E2 ;
                        10'h37A : QQ <= 9'h0E1 ;
                        10'h37B : QQ <= 9'h0E0 ;
                        10'h37C : QQ <= 9'h0DE ;
                        10'h37D : QQ <= 9'h0DD ;
                        10'h37E : QQ <= 9'h0DB ;
                        10'h37F : QQ <= 9'h0DA ;
                        10'h380 : QQ <= 9'h0D9 ;
                        10'h381 : QQ <= 9'h0D7 ;
                        10'h382 : QQ <= 9'h0D6 ;
                        10'h383 : QQ <= 9'h0D4 ;
                        10'h384 : QQ <= 9'h0D3 ;
                        10'h385 : QQ <= 9'h0D2 ;
                        10'h386 : QQ <= 9'h0D0 ;
                        10'h387 : QQ <= 9'h0CF ;
                        10'h388 : QQ <= 9'h0CD ;
                        10'h389 : QQ <= 9'h0CC ;
                        10'h38A : QQ <= 9'h0CB ;
                        10'h38B : QQ <= 9'h0C9 ;
                        10'h38C : QQ <= 9'h0C8 ;
                        10'h38D : QQ <= 9'h0C6 ;
                        10'h38E : QQ <= 9'h0C5 ;
                        10'h38F : QQ <= 9'h0C3 ;
                        10'h390 : QQ <= 9'h0C2 ;
                        10'h391 : QQ <= 9'h0C0 ;
                        10'h392 : QQ <= 9'h0BF ;
                        10'h393 : QQ <= 9'h0BD ;
                        10'h394 : QQ <= 9'h0BC ;
                        10'h395 : QQ <= 9'h0BA ;
                        10'h396 : QQ <= 9'h0B9 ;
                        10'h397 : QQ <= 9'h0B7 ;
                        10'h398 : QQ <= 9'h0B6 ;
                        10'h399 : QQ <= 9'h0B4 ;
                        10'h39A : QQ <= 9'h0B3 ;
                        10'h39B : QQ <= 9'h0B1 ;
                        10'h39C : QQ <= 9'h0B0 ;
                        10'h39D : QQ <= 9'h0AE ;
                        10'h39E : QQ <= 9'h0AD ;
                        10'h39F : QQ <= 9'h0AB ;
                        10'h3A0 : QQ <= 9'h0AA ;
                        10'h3A1 : QQ <= 9'h0A8 ;
                        10'h3A2 : QQ <= 9'h0A7 ;
                        10'h3A3 : QQ <= 9'h0A5 ;
                        10'h3A4 : QQ <= 9'h0A4 ;
                        10'h3A5 : QQ <= 9'h0A2 ;
                        10'h3A6 : QQ <= 9'h0A1 ;
                        10'h3A7 : QQ <= 9'h09F ;
                        10'h3A8 : QQ <= 9'h09D ;
                        10'h3A9 : QQ <= 9'h09C ;
                        10'h3AA : QQ <= 9'h09A ;
                        10'h3AB : QQ <= 9'h099 ;
                        10'h3AC : QQ <= 9'h097 ;
                        10'h3AD : QQ <= 9'h095 ;
                        10'h3AE : QQ <= 9'h094 ;
                        10'h3AF : QQ <= 9'h092 ;
                        10'h3B0 : QQ <= 9'h091 ;
                        10'h3B1 : QQ <= 9'h08F ;
                        10'h3B2 : QQ <= 9'h08D ;
                        10'h3B3 : QQ <= 9'h08C ;
                        10'h3B4 : QQ <= 9'h08A ;
                        10'h3B5 : QQ <= 9'h088 ;
                        10'h3B6 : QQ <= 9'h087 ;
                        10'h3B7 : QQ <= 9'h085 ;
                        10'h3B8 : QQ <= 9'h084 ;
                        10'h3B9 : QQ <= 9'h082 ;
                        10'h3BA : QQ <= 9'h080 ;
                        10'h3BB : QQ <= 9'h07F ;
                        10'h3BC : QQ <= 9'h07D ;
                        10'h3BD : QQ <= 9'h07B ;
                        10'h3BE : QQ <= 9'h07A ;
                        10'h3BF : QQ <= 9'h078 ;
                        10'h3C0 : QQ <= 9'h076 ;
                        10'h3C1 : QQ <= 9'h074 ;
                        10'h3C2 : QQ <= 9'h073 ;
                        10'h3C3 : QQ <= 9'h071 ;
                        10'h3C4 : QQ <= 9'h06F ;
                        10'h3C5 : QQ <= 9'h06E ;
                        10'h3C6 : QQ <= 9'h06C ;
                        10'h3C7 : QQ <= 9'h06A ;
                        10'h3C8 : QQ <= 9'h068 ;
                        10'h3C9 : QQ <= 9'h067 ;
                        10'h3CA : QQ <= 9'h065 ;
                        10'h3CB : QQ <= 9'h063 ;
                        10'h3CC : QQ <= 9'h061 ;
                        10'h3CD : QQ <= 9'h060 ;
                        10'h3CE : QQ <= 9'h05E ;
                        10'h3CF : QQ <= 9'h05C ;
                        10'h3D0 : QQ <= 9'h05A ;
                        10'h3D1 : QQ <= 9'h059 ;
                        10'h3D2 : QQ <= 9'h057 ;
                        10'h3D3 : QQ <= 9'h055 ;
                        10'h3D4 : QQ <= 9'h053 ;
                        10'h3D5 : QQ <= 9'h052 ;
                        10'h3D6 : QQ <= 9'h050 ;
                        10'h3D7 : QQ <= 9'h04E ;
                        10'h3D8 : QQ <= 9'h04C ;
                        10'h3D9 : QQ <= 9'h04A ;
                        10'h3DA : QQ <= 9'h049 ;
                        10'h3DB : QQ <= 9'h047 ;
                        10'h3DC : QQ <= 9'h045 ;
                        10'h3DD : QQ <= 9'h043 ;
                        10'h3DE : QQ <= 9'h041 ;
                        10'h3DF : QQ <= 9'h03F ;
                        10'h3E0 : QQ <= 9'h03E ;
                        10'h3E1 : QQ <= 9'h03C ;
                        10'h3E2 : QQ <= 9'h03A ;
                        10'h3E3 : QQ <= 9'h038 ;
                        10'h3E4 : QQ <= 9'h036 ;
                        10'h3E5 : QQ <= 9'h034 ;
                        10'h3E6 : QQ <= 9'h032 ;
                        10'h3E7 : QQ <= 9'h030 ;
                        10'h3E8 : QQ <= 9'h02F ;
                        10'h3E9 : QQ <= 9'h02D ;
                        10'h3EA : QQ <= 9'h02B ;
                        10'h3EB : QQ <= 9'h029 ;
                        10'h3EC : QQ <= 9'h027 ;
                        10'h3ED : QQ <= 9'h025 ;
                        10'h3EE : QQ <= 9'h023 ;
                        10'h3EF : QQ <= 9'h021 ;
                        10'h3F0 : QQ <= 9'h01F ;
                        10'h3F1 : QQ <= 9'h01D ;
                        10'h3F2 : QQ <= 9'h01C ;
                        10'h3F3 : QQ <= 9'h01A ;
                        10'h3F4 : QQ <= 9'h018 ;
                        10'h3F5 : QQ <= 9'h016 ;
                        10'h3F6 : QQ <= 9'h014 ;
                        10'h3F7 : QQ <= 9'h012 ;
                        10'h3F8 : QQ <= 9'h010 ;
                        10'h3F9 : QQ <= 9'h00E ;
                        10'h3FA : QQ <= 9'h00C ;
                        10'h3FB : QQ <= 9'h00A ;
                        10'h3FC : QQ <= 9'h008 ;
                        10'h3FD : QQ <= 9'h006 ;
                        10'h3FE : QQ <= 9'h004 ;
                        10'h3FF : QQ <= 9'h002 ;
                endcase
        assign QQ_o = QQ ;
endmodule // SIN_ROM_4s11_s11

